module bus(

);

reg bus[0:7];



